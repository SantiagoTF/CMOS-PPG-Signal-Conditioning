** sch_path: /home/designer/shared/Design/CCLNA/testbench_CurrentM_OTA.sch
**.subckt testbench_CurrentM_OTA
XM3 net5 net1 VDD VDD sg13_hv_pmos w=4u l=1u ng=1 m=3
XM5 net2 net2 VDD VDD sg13_hv_pmos w=4u l=1u ng=1 m=1
XM6 VOut net2 VDD VDD sg13_hv_pmos w=4u l=1u ng=1 m=3
XM7 net1 Vin- net3 net3 sg13_hv_nmos w=8u l=1u ng=1 m=1
XM8 net2 Vin+ net3 net3 sg13_hv_nmos w=8u l=1u ng=1 m=1
XM9 net3 net4 VSS VSS sg13_hv_nmos w=2u l=1u ng=1 m=1
XM10 net4 net4 VSS VSS sg13_hv_nmos w=2u l=1u ng=1 m=1
XM11 net5 net5 VSS VSS sg13_hv_nmos w=3u l=1u ng=1 m=1
XM12 VOut net5 VSS VSS sg13_hv_nmos w=3u l=1u ng=1 m=1
I0 VDD net4 2u
E1 Vin- net7 net6 VSS -0.5
E2 Vin+ net7 net6 VSS 0.5
V1 net7 GND 0.4
V2 net6 GND dc 0 ac 1 sin(0 8m 100k)
V3 VDD GND 3.3
V4 VSS GND 0
C1 VOut VSS 5p m=1
XM4 net1 net1 VDD VDD sg13_hv_pmos w=4u l=1u ng=1 m=1
**** begin user architecture code
 .lib cornerMOShv.lib mos_tt


.param temp=27
.save all

.control
  ac dec 80 0.1 11g
  set filetype = ascii
  set units=degrees
  write testbench_CurrentM_OTA.raw vdb(vout) vp(vout)
  set appendwrite
  op
  set filetype = ascii
  write testbench_CurrentM_OTA.raw

  * tran 0.1u 100u
  * set filetype = ascii
  * write testbench_CurrentM_OTA.raw v(vin+) v(vin-) v(vout)
  * set appendwrite
  * op
  * set filetype = ascii
  * write testbench_CurrentM_OTA.raw

.endc


**** end user architecture code
**.ends
.GLOBAL GND
.end
